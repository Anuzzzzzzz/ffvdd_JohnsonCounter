`include "transaction.sv"
`include "generator.sv"
`include "bfm.sv"
`include "interface.sv"
`include "environment.sv"
`include "test.sv"
`include "design.v"
`include "assert_jc.sv"
`include "testbench.sv"
