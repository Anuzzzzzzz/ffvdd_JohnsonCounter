class transaction;
bit [7:0] q;
function void display();
$display("------------------------------------------------------------------------ ");
$display(" \t q= %0b",q);
$display(" ------------------------------------------------------------------------");

endfunction
endclass
